`define RV64
`define RV_PMU_PORTS
`define RV_SCAN_PORTS
`define RV_TRACE_PORTS
`define RV_BUILD_ETRACE
`define RV_ICACHE_MAX_ENTRIES 1024
`define RV_ICACHE_ENABLE
`define RV_DC_ENABLE
`define RV_DCPREF_ENABLE
`define RV_DC_NUM_BANKS 16
`define RV_NO_SECONDARY_ALU
`define RV_BUILD_FPU
`define RV_BUILD_BITMANIP
`define RV_DATA_GATING
`define RV_AXI_BUS_DATAWIDTH 512
`define OOO_ENABLE
`define RV_OOO_ISSQ_DEPTH 17
`define RV_OOO_STISSQ_DEPTH 24
`define RV_OOO_CHKPTTOTAL 24
`define RV_BHT_SIZE 2048
`define RV_BTB_SIZE 512
`define RV_BTB_WAYS 4
`define RV_BTB_BTAG_SIZE_LIMIT 22
`define RV_BROFFSET_WIDTH 20
`define RV_BTB2_ENABLE
`define RV_BTB2_ARRAY_DEPTH 128
`define RV_BTB2_WAYS 3
`define NPC_ENABLE
`define NPC_ENTRIES 16
`define NPC_INDEX_MODE
`define NPC2_ENTRIES 128
`define ALN_xFB_SIZE 1
`define TAGE_ENABLE
`define TAGE_TABLES 5
`define TAGE_ENTRIES 2048
`define TAGE_RAM_ENABLE
`define TAGE_CACHE_WAY 5
`define TAGE_CACHE_ENTRIES 256
`define TAGE_CACHE_GFOLD_TABLE_IDX 2
`define BIG_TAGE_NUM_BANKS_PER_TABLE 4
`define BIG_TAGE_NUM_WAYS 2
`define RV_BTBI_ENABLE
`define RV_BTBI_CONST_ENABLE
`define RV_CCB_ENABLE
`define RAS_ENABLE
`define RV_BUILD_VEU
`define RV_VEU_MAX_VL 128
`define RV_PRIVATE_L2
`define RV_PL2_SIZE 256
`define PL2_TAG_BANKING_ENABLE
`define RV_L2_PREF_ENABLE
`define L2PREF_RST_STRIDE_DEGREE 4
`define RV_PL2_PB_DEPTH 32
`define RV_PL2_ECC_ENABLE
`define IFU_PL2_ACCESS_EN
`define ITLB_NUM_ENTRIES 64
`define RV_BUILD_VCRYPTO
`define AXI_ASYNC_OUTPUTS
`define RV_BUILD_HYPERVISOR
`define RV_NUM_PMP 16
`define RV_BUILD_KRYPTO
`define RV_AXI_BUS_TAG 7
`define RV_LSU_NUM_NBLOAD 16
`define PW_CACHE_ENABLE
`define RV_LDST_PER_CYCLE 3
`define RV_LD_PER_CYCLE 2
`define ITTAGE_ENABLE
`define RV_ICACHE_SIZE 64
`define RV_DC_SIZE 64
`define RV_INST_FETCH_WIDTH 16
`define RV_DEC_INSTBUF_DEPTH 16
`define RV_DEC_DISPATCH_WIDTH 6
`define RV_DEC_DISPATCH_PIPESTAGE_DP2_ENABLE
`define RV_ALN_DEC_USECREDITS
`define RV_OOO_NUM_ALU_ISSQ 6
`define RV_OOO_LRQD 75
`define RV_OOO_NPR 192
`define RV_OOO_ROBD 259
`define RV_OOO_SRQD 66
`define RV_OOO_VLIQD 32
`define RV_OOO_VSIQD 24
`define DTLB_NUM_ENTRIES 64
`define DTLB_SAM_DEC
`define MMU_SIZE 2048
`define RV_DCPREF_OOO_LIMIT 64
`define RV_DCPREF_PRQSIZE 64
`define RV_BUILD_AIA_WIREDONLY
`define RV_BUILD_REAL_TIME
`define RV_BUILD_SSTC
`define CORESIGHT_ENABLE
`define RV_IO_ATOMIC
`define STRUCTURAL_GPR_ENABLE
`define ACLINT_EXT_OR_INT
`define ASSERT_ON
`define AXI_ASYNC_FIFO_STORE SRAM
`define BIG_TAGE
`define BIG_TAGE_10_TWOWAY 0
`define BIG_TAGE_11_TWOWAY 0
`define BIG_TAGE_12_TWOWAY 0
`define BIG_TAGE_13_TWOWAY 0
`define BIG_TAGE_14_TWOWAY 0
`define BIG_TAGE_1_TWOWAY 0
`define BIG_TAGE_2_TWOWAY 0
`define BIG_TAGE_3_TWOWAY 0
`define BIG_TAGE_4_TWOWAY 0
`define BIG_TAGE_5_TWOWAY 0
`define BIG_TAGE_6_TWOWAY 0
`define BIG_TAGE_7_TWOWAY 0
`define BIG_TAGE_8_TWOWAY 0
`define BIG_TAGE_9_TWOWAY 0
`define CACHE_LINE_SIZE 64
`define CCB_NUM_NCWR_PERSRC 2
`define CLOCK_PERIOD 100
`define CPU_TOP `RV_TOP.shasta
`define CS_ARCH_CODE 32'hdc100000
`define CS_AUTHSTATUS 13'hfb8
`define CS_CIDR0 13'hff0
`define CS_CIDR1 13'hff4
`define CS_CIDR2 13'hff8
`define CS_CIDR3 13'hffc
`define CS_CLAIMCLR 13'hfa4
`define CS_CLAIMSET 13'hfa0
`define CS_COMP_CLASS 4'he
`define CS_COMP_ID0 32'hd
`define CS_COMP_ID2 32'h5
`define CS_COMP_ID3 32'hb1
`define CS_DESIGN_REV 4'h0
`define CS_DEVAFF0 13'hfa8
`define CS_DEVAFF1 13'hfac
`define CS_DEVARCH 13'hfbc
`define CS_DEVICE_AFF0 32'h0
`define CS_DEVICE_AFF1 32'h0
`define CS_DEVICE_ID 32'h0
`define CS_DEVICE_ID1 32'h0
`define CS_DEVICE_ID2 32'h0
`define CS_DEVICE_PN 12'h0
`define CS_DEVID 13'hfc8
`define CS_DEVID1 13'hfc4
`define CS_DEVID2 13'hfc0
`define CS_DEVTYPE 13'hfcc
`define CS_ERRATA_REV 4'h0
`define CS_ITCTRL 13'hf00
`define CS_LAR 13'hfb0
`define CS_LSR 13'hfb4
`define CS_MOD_REV 4'h0
`define CS_PERIPH_ID5 32'h0
`define CS_PERIPH_ID6 32'h0
`define CS_PERIPH_ID7 32'h0
`define CS_PIDR0 13'hfe0
`define CS_PIDR1 13'hfe4
`define CS_PIDR2 13'hfe8
`define CS_PIDR3 13'hfec
`define CS_PIDR4 13'hfd0
`define CS_PIDR5 13'hfd4
`define CS_PIDR6 13'hfd8
`define CS_PIDR7 13'hfdc
`define CS_TYPE_DEBUG 4'h5
`define CS_TYPE_PROC 4'h1
`define DATAWIDTH 64
`define DEC_ASSERT
`define DTLB_NUM_ENTRIES_FINAL 64
`define DTLB_NUM_SETS_1G 2
`define DTLB_NUM_SETS_2M 8
`define DTLB_NUM_SETS_4K 16
`define DTLB_NUM_WAYS 4
`define DTLB_SAM_DEC_ENABLE
`define DTLB_SET_ENABLE
`define EXU_SLOTS_WIDTH 6
`define FPU_ASSERT2COV
`define FPU_EXTERNAL_FPR
`define GPA_SIZE 59
`define GPA_VPN_SIZE 47
`define IC_NUM_WAYS 4
`define IC_ROW_INC 0
`define IFU_AXI_WIDTH_512 1
`define IFU_AXI_WIDTH_NEQ_64 1
`define ITLB_NUM_SETS_1G 2
`define ITLB_NUM_SETS_2M 8
`define ITLB_NUM_SETS_4K 16
`define ITLB_NUM_WAYS 4
`define ITLB_SET_ENABLE
`define ITTAGE_ENTRIES 512
`define ITTAGE_ENTRY_INDEX 9
`define ITTAGE_HIST_0 2
`define ITTAGE_HIST_1 16
`define ITTAGE_HIST_2 128
`define ITTAGE_RTL_ENABLE
`define ITTAGE_TABLES 3
`define ITTAGE_TAG_WIDTH 12
`define ITTAGE_U_ALLOC_SET_ENABLE
`define ITTAGE_U_WIDTH 2
`define L2PREF_FIFO_DEPTH 16
`define L2PREF_NUM_ENT 64
`define L2PREF_NUM_STRIDES 4
`define L2PREF_RST_PAGE_XING 0
`define L2PREF_STRIDE_SIZE 12
`define L2PREF_TAG_SIZE 12
`define L2PREF_WAYS 4
`define LSU_AXI_WIDTH_512 1
`define LSU_BUSW_EQ_CLW 1
`define MAILBOX_ADDR 64'hd0580000
`define MMU_ASID_ARRAY_SIZE 30
`define MMU_ENABLE
`define MMU_ENTRIES 512
`define MMU_GPA_ARRAY_SIZE 70
`define MMU_HFENCE_OPTIMIZATION
`define MMU_IFU_PWQ_ENTRIES 4
`define MMU_IFU_PWQ_PTR_BITS 2
`define MMU_INDEX_BITS 9
`define MMU_LSU_PWQ_ENTRIES 4
`define MMU_LSU_PWQ_PTR_BITS 2
`define MMU_NUM_IFU_PW_1
`define MMU_NUM_LSU_PW_2
`define MMU_NUM_PAGEWALKS 3
`define MMU_NUM_PAGEWALKS_IFU 1
`define MMU_NUM_PAGEWALKS_IFU_FINAL 1
`define MMU_NUM_PAGEWALKS_LSU 2
`define MMU_NUM_PAGEWALKS_LSU_FINAL 2
`define MMU_NUM_PROPS 18
`define MMU_PAGESIZES 5
`define MMU_PWQ_ENABLE
`define MMU_TAG_PROPS 7
`define MMU_TAG_SIZE 50
`define MMU_WAYS 4
`define NPC_CONF_INST_VAL 3
`define NPC_CONF_WIDTH 2
`define NPC_ENABLE_FINAL
`define NPC_TAG_WIDTH 12
`define NPC_TGT_WIDTH 12
`define NPC_USE_INST_VAL 1
`define NUM_CORES 1
`define NUM_CORES_1
`define NUM_HARTS 1
`define NUM_THREADS 1
`define NUM_THREADS_LOG 0
`define PA_ALL_ZEROES 39'h0
`define PA_MASK 39'h7fffffffff
`define PA_SIZE 39
`define PL2_DC_NBANKS 2
`define PROGBUF_NUM 0
`define PWC_ENABLE
`define PWC_ENTRIES 32
`define RAS_CNT_INC_DEC
`define RAS_DEPTH 128
`define RAS_INDEX 7
`define RAS_OOO_ENABLE
`define REAL_COMM_ENABLE
`define REAL_COMM_RS
`define RV32_CLINT_BASE_ADDR 34'hdc001000
`define RV32_PLIC_BASE_ADDR 34'hd8000000
`define RV32_PLIC_IP_BASE_ADDR 34'hdc000000
`define RV64_CLINT_BASE_ADDR 64'h68dc001000
`define RV64_PLIC_BASE_ADDR 64'h68d8000000
`define RV64_PLIC_IP_BASE_ADDR 64'h68dc000000
`define RV64_VA57
`define RV_ADD_ADDL_FLOP
`define RV_AIA_IMSIC_INT_FILE_BASE_OFFSET 19'h0
`define RV_AIA_IMSIC_MFILE_BASE_ADDR 39'h0
`define RV_AIA_IMSIC_MFILE_SIZE 4
`define RV_AIA_IMSIC_SFILE_BASE_ADDR 39'h0
`define RV_AIA_IMSIC_SFILE_SIZE 4
`define RV_AIA_MSI_NUM_INTERRUPT_IDS 63
`define RV_AIA_NONIMSIC_CSRS_EXIST
`define RV_AMU_BUF_DEPTH 1024
`define RV_AMU_EVENTS_NUM 43
`define RV_AMU_SADR 23'h441000
`define RV_AMU_SIZE 256
`define RV_AXI_ONE_BEAT_RETURN
`define RV_AXI_SIZE_WIDTH 3
`define RV_BHT_ADDR_HI 11
`define RV_BHT_ADDR_LO 5
`define RV_BHT_ARRAY_DEPTH 128
`define RV_BHT_GHR_PAD fghr[123:0],3'b0
`define RV_BHT_GHR_PAD2 fghr[124:0],2'b0
`define RV_BHT_GHR_RANGE 127:0
`define RV_BHT_GHR_SIZE 128
`define RV_BHT_HASH_STRING {ghr[126:6] ^ {ghr[126+1], {127-1-6{1'b0} } },hashin[9:4]^ghr[6-1:0]}
`define RV_BHT_NUM_BANKS 16
`define RV_BHT_SIZE_LOG 11
`define RV_BP_FETCH_WIDTH 16
`define RV_BTB2_ADDR_HI 11
`define RV_BTB2_ADDR_LO 5
`define RV_BTB2_BTAG_FOLD 1
`define RV_BTB2_BTAG_SIZE 14
`define RV_BTB2_BTAG_SIZE_LIMIT 22
`define RV_BTB2_DATA_SIZE 41
`define RV_BTB2_DPRAM_ENABLE
`define RV_BTB2_DPRAM_SIZE 8192
`define RV_BTB2_INDEX1_HI 11
`define RV_BTB2_INDEX1_LO 5
`define RV_BTB2_SIZE 2048
`define RV_BTBI_ADDR_HI 13
`define RV_BTBI_ADDR_LO 5
`define RV_BTBI_ARRAY_DEPTH 512
`define RV_BTBI_CONST_ADDR_HI 12
`define RV_BTBI_CONST_ADDR_LO 5
`define RV_BTBI_CONST_SIZE 256
`define RV_BTBI_CONST_TAG_SIZE 13
`define RV_BTBI_CONST_WAYS 2
`define RV_BTBI_DATA_SIZE 63
`define RV_BTBI_SIZE 512
`define RV_BTB_ADDR_HI 9
`define RV_BTB_ADDR_LO 5
`define RV_BTB_ARRAY_DEPTH 32
`define RV_BTB_BTAG_SIZE 13
`define RV_BTB_DATA_SIZE 40
`define RV_BTB_INDEX1_HI 9
`define RV_BTB_INDEX1_LO 5
`define RV_BTB_INDEX2_HI 15
`define RV_BTB_INDEX2_LO 10
`define RV_BTB_INDEX3_HI 21
`define RV_BTB_INDEX3_LO 16
`define RV_BUILD_AFFINITY_REGISTER
`define RV_BUILD_AIA
`define RV_BUILD_AMO
`define RV_BUILD_AXI4 1
`define RV_BUILD_ETRACEorRV_TRACE_PORTS
`define RV_BUILD_EXTINT_PORTS
`define RV_BUILD_EXT_TIMER
`define RV_BUILD_FPU_BF16
`define RV_BUILD_FPU_FP16
`define RV_BUILD_FPU_ZFA
`define RV_BUILD_KRYPTO_BIT
`define RV_BUILD_KRYPTO_NIST
`define RV_BUILD_KRYPTO_SM
`define RV_BUILD_SWINT
`define RV_BUILD_VCRYPTO_BIT
`define RV_BUILD_VCRYPTO_NIST
`define RV_BUILD_VCRYPTO_SM
`define RV_BUILD_ZABHA
`define RV_BUILD_ZACAS
`define RV_BUILD_ZBA
`define RV_BUILD_ZBB
`define RV_BUILD_ZBC
`define RV_BUILD_ZBKB
`define RV_BUILD_ZBKC
`define RV_BUILD_ZBKX
`define RV_BUILD_ZBS
`define RV_BUILD_ZCB
`define RV_BUILD_ZICOND
`define RV_BUILD_ZK
`define RV_BUILD_ZKND
`define RV_BUILD_ZKNE
`define RV_BUILD_ZKNED
`define RV_BUILD_ZKNH
`define RV_BUILD_ZKSED
`define RV_BUILD_ZKSH
`define RV_BUILD_ZVBB
`define RV_BUILD_ZVBC
`define RV_BUILD_ZVKB
`define RV_BUILD_ZVKG
`define RV_BUILD_ZVKNED
`define RV_BUILD_ZVKNHA
`define RV_BUILD_ZVKNHB
`define RV_BUILD_ZVKSED
`define RV_BUILD_ZVKSH
`define RV_BUS_BYTEWIDTH 64
`define RV_CLINT_BASE_ADDR 39'h68dc001000
`define RV_CLINT_SIZE 39'h10f00
`define RV_CONFIGPTR 39'h0
`define RV_DATA_ACCESS_ADDR0 39'h0
`define RV_DATA_ACCESS_ADDR1 39'h0
`define RV_DATA_ACCESS_ADDR2 39'h0
`define RV_DATA_ACCESS_ADDR3 39'h0
`define RV_DATA_ACCESS_ADDR4 39'h0
`define RV_DATA_ACCESS_ADDR5 39'h0
`define RV_DATA_ACCESS_ADDR6 39'h0
`define RV_DATA_ACCESS_ADDR7 39'h0
`define RV_DATA_ACCESS_ENABLE0 1'h0
`define RV_DATA_ACCESS_ENABLE1 1'h0
`define RV_DATA_ACCESS_ENABLE2 1'h0
`define RV_DATA_ACCESS_ENABLE3 1'h0
`define RV_DATA_ACCESS_ENABLE4 1'h0
`define RV_DATA_ACCESS_ENABLE5 1'h0
`define RV_DATA_ACCESS_ENABLE6 1'h0
`define RV_DATA_ACCESS_ENABLE7 1'h0
`define RV_DATA_ACCESS_MASK0 39'h7fffffffff
`define RV_DATA_ACCESS_MASK1 39'h7fffffffff
`define RV_DATA_ACCESS_MASK2 39'h7fffffffff
`define RV_DATA_ACCESS_MASK3 39'h7fffffffff
`define RV_DATA_ACCESS_MASK4 39'h7fffffffff
`define RV_DATA_ACCESS_MASK5 39'h7fffffffff
`define RV_DATA_ACCESS_MASK6 39'h7fffffffff
`define RV_DATA_ACCESS_MASK7 39'h7fffffffff
`define RV_DATA_GATING_LOW_FREQ_WIDTH 4
`define RV_DBG_VER1P0
`define RV_DCACHE_LINE_SIZE 64
`define RV_DCCM_ARRAY_SIZE 2
`define RV_DCCM_BANK_BITS 5
`define RV_DCCM_BITS 16
`define RV_DCCM_BYTE_WIDTH 4
`define RV_DCCM_DATA_CELL ram_512x39
`define RV_DCCM_DATA_WIDTH 32
`define RV_DCCM_EADR 39'h780004ffff
`define RV_DCCM_ECC_ENABLE
`define RV_DCCM_ECC_WIDTH 7
`define RV_DCCM_FDATA_WIDTH 39
`define RV_DCCM_HI_ARRAY_SIZE 1
`define RV_DCCM_HI_BANK_BITS 0
`define RV_DCCM_HI_DATA_CELL ram_256x39
`define RV_DCCM_HI_INDEX_BITS 8
`define RV_DCCM_HI_ROWS 256
`define RV_DCCM_INDEX_BITS 9
`define RV_DCCM_LO_ARRAY_SIZE 2
`define RV_DCCM_LO_BANK_BITS 2
`define RV_DCCM_LO_DATA_CELL ram_512x39
`define RV_DCCM_LO_INDEX_BITS 9
`define RV_DCCM_LO_ROWS 512
`define RV_DCCM_NUM_BANKS 32
`define RV_DCCM_NUM_BANKS_32
`define RV_DCCM_NUM_HI_BANKS 1
`define RV_DCCM_NUM_LO_BANKS 4
`define RV_DCCM_OFFSET 28'h40000
`define RV_DCCM_REGION 4'hf
`define RV_DCCM_RESERVED 'h1000
`define RV_DCCM_ROWS 512
`define RV_DCCM_SADR 39'h7800040000
`define RV_DCCM_SEL_HI_BANKS 0
`define RV_DCCM_SIZE 64
`define RV_DCCM_SIZE_64
`define RV_DCCM_SIZE_NON_POWER_TWO 0
`define RV_DCCM_SIZE_NON_POWER_TWO_0
`define RV_DCCM_WIDTH_BITS 2
`define RV_DC_DATA_CELL ram_1024x39
`define RV_DC_NUM_ROWS 1024
`define RV_DC_NUM_WAYS 16
`define RV_DEBUG_SB_MEM 'hb0580000
`define RV_DEC_DISPATCH_WIDTH_GREATER_EQUAL_2
`define RV_DEC_DISPATCH_WIDTH_GREATER_EQUAL_3
`define RV_DEC_DISPATCH_WIDTH_GREATER_EQUAL_4
`define RV_DMA_BUF_DEPTH 4
`define RV_DMA_BUS_TAG 1
`define RV_EXTERNAL_DATA 'hc0580000
`define RV_EXTERNAL_DATA_1 'h0
`define RV_EXTERNAL_PROG 'hb0000000
`define RV_EXT_ADDRWIDTH 32
`define RV_EXT_DATAWIDTH 64
`define RV_GEILEN 0
`define RV_HARTID_WIDTH 8
`define RV_HASH_LT_DELTA
`define RV_HASH_LT_GHR
`define RV_ICACHE_DATA_CELL ram_512x34
`define RV_ICACHE_IC_DEPTH 10
`define RV_ICACHE_IC_INDEX 10
`define RV_ICACHE_IC_ROWS 512
`define RV_ICACHE_LINE_SIZE 64
`define RV_ICACHE_TADDR_HIGH 7
`define RV_ICACHE_TAG_CELL ram_256x28
`define RV_ICACHE_TAG_DEPTH 256
`define RV_ICACHE_TAG_HIGH 14
`define RV_ICACHE_TAG_LOW 6
`define RV_ICACHE_TAG_WIDTH 28
`define RV_ICACHE_WDATA_WIDTH 272
`define RV_ICCM_2_LVL_MUX_ENABLE
`define RV_ICCM_BANK_BITS 8
`define RV_ICCM_BITS 19
`define RV_ICCM_DATA_CELL ram_512x39
`define RV_ICCM_EADR 39'h700e07ffff
`define RV_ICCM_ECC
`define RV_ICCM_HI_BANKS_DATA_CELL ram_0x39
`define RV_ICCM_HI_BANKS_INDEX_BITS 0
`define RV_ICCM_HI_BANKS_MACRO_ENTRIES 0
`define RV_ICCM_HI_BANKS_MACRO_SIZE 0
`define RV_ICCM_HI_BANKS_SIZE 0
`define RV_ICCM_INDEX_BITS 9
`define RV_ICCM_INDEX_BITS_PRELIM 15
`define RV_ICCM_MAX_INDEX_BITS 9
`define RV_ICCM_MAX_MACRO_ENTRIES 512
`define RV_ICCM_MAX_MACRO_SIZE 2
`define RV_ICCM_MIN_X_BANKS 2
`define RV_ICCM_NON_POWER_TWO_SIZE_512_512
`define RV_ICCM_NUM_BANKS 256
`define RV_ICCM_NUM_BANKS_256
`define RV_ICCM_NUM_Y_BANKS 64
`define RV_ICCM_NUM_Y_BANKS_LO 64
`define RV_ICCM_OFFSET 10'he000000
`define RV_ICCM_REGION 4'he
`define RV_ICCM_RESERVED 'h1000
`define RV_ICCM_ROWS 512
`define RV_ICCM_SADR 39'h700e000000
`define RV_ICCM_SIZE 512
`define RV_ICCM_SIZE_512
`define RV_IC_BLOCKS 1
`define RV_IFUFW_IS_16
`define RV_IFU_BUS_DATAWIDTH 512
`define RV_IFU_BUS_TAG 3
`define RV_IFU_MB_ENTRIES 8
`define RV_IFU_PREFETCH_ENABLE
`define RV_INDIR_CSRS_EXIST
`define RV_INST_ACCESS_ADDR0 39'h0
`define RV_INST_ACCESS_ADDR1 39'h0
`define RV_INST_ACCESS_ADDR2 39'h0
`define RV_INST_ACCESS_ADDR3 39'h0
`define RV_INST_ACCESS_ADDR4 39'h0
`define RV_INST_ACCESS_ADDR5 39'h0
`define RV_INST_ACCESS_ADDR6 39'h0
`define RV_INST_ACCESS_ADDR7 39'h0
`define RV_INST_ACCESS_ENABLE0 1'h0
`define RV_INST_ACCESS_ENABLE1 1'h0
`define RV_INST_ACCESS_ENABLE2 1'h0
`define RV_INST_ACCESS_ENABLE3 1'h0
`define RV_INST_ACCESS_ENABLE4 1'h0
`define RV_INST_ACCESS_ENABLE5 1'h0
`define RV_INST_ACCESS_ENABLE6 1'h0
`define RV_INST_ACCESS_ENABLE7 1'h0
`define RV_INST_ACCESS_MASK0 39'h7fffffffff
`define RV_INST_ACCESS_MASK1 39'h7fffffffff
`define RV_INST_ACCESS_MASK2 39'h7fffffffff
`define RV_INST_ACCESS_MASK3 39'h7fffffffff
`define RV_INST_ACCESS_MASK4 39'h7fffffffff
`define RV_INST_ACCESS_MASK5 39'h7fffffffff
`define RV_INST_ACCESS_MASK6 39'h7fffffffff
`define RV_INST_ACCESS_MASK7 39'h7fffffffff
`define RV_IOF_EADR 39'h2800000fff
`define RV_IOF_SADR 39'h2800000000
`define RV_IOF_SIZE 4
`define RV_ITS_EADR 39'h7800003fff
`define RV_ITS_REG_EADR 39'h4000003fff
`define RV_ITS_REG_SADR 39'h4000000000
`define RV_ITS_REG_SIZE 16
`define RV_ITS_SADR 39'h7800000000
`define RV_ITS_SIZE 16
`define RV_LDERR_ROLLBACK 1
`define RV_LSU_BUS_DATAWIDTH 512
`define RV_LSU_BUS_TAG 7
`define RV_LSU_DATA_WIDTH 128
`define RV_LSU_ECC_ENABLE
`define RV_LSU_NUM_NBLOAD_WIDTH 4
`define RV_LSU_SB_BITS 16
`define RV_LSU_STBUF_DEPTH 8
`define RV_MISALIGN_ENABLE
`define RV_MPC_PORTS
`define RV_MSIP_BASE_ADDR 39'h78000d8000
`define RV_MSIP_BITS 14
`define RV_MSIP_OFFSET 'hd8000
`define RV_MSIP_REGION 'hf
`define RV_MSIP_SIZE 16
`define RV_MSI_LAST_INTERRUPT_ID_FOR_PCIE 2047
`define RV_MSI_STARTING_INTERRUPT_ID_FOR_PCIE 1024
`define RV_MTIMECMP_BASE_ADDR 39'h78000d0000
`define RV_MTIMECMP_BITS 15
`define RV_MTIMECMP_OFFSET 'hd0000
`define RV_MTIMECMP_REGION 'hf
`define RV_MTIMECMP_SIZE 32
`define RV_MTIMER_BASE_ADDR 39'h78000c8000
`define RV_MTIMER_BITS 15
`define RV_MTIMER_OFFSET 'hc8000
`define RV_MTIMER_REGION 'hf
`define RV_MTIMER_SIZE 32
`define RV_MULTIPLE_LDST_PER_CYCLE
`define RV_MVENDORID_BANK 13
`define RV_MVENDORID_OFFSET 96
`define RV_NHPM 4
`define RV_NMI_VEC 39'hee000000
`define RV_NUMIREGS 32
`define RV_NUM_STATEEN 4
`define RV_OOO_CHKPTPERCYC 2
`define RV_OOO_FVNPR 128
`define RV_OOO_INPR 192
`define RV_OOO_NPRVS 32
`define RV_OOO_NUM_FPU_ISSQ 2
`define RV_OOO_NUM_VEU_ISSQ 2
`define RV_PD_PARTITION
`define RV_PIC_BASE_ADDR 39'h78000c0000
`define RV_PIC_BITS 15
`define RV_PIC_INT_WORDS 1
`define RV_PIC_MEIE_COUNT 12
`define RV_PIC_MEIE_MASK 'h1
`define RV_PIC_MEIE_OFFSET 'h2000
`define RV_PIC_MEIGWCLR_COUNT 12
`define RV_PIC_MEIGWCLR_MASK 'h0
`define RV_PIC_MEIGWCLR_OFFSET 'h5000
`define RV_PIC_MEIGWCTRL_COUNT 12
`define RV_PIC_MEIGWCTRL_MASK 'h3
`define RV_PIC_MEIGWCTRL_OFFSET 'h4000
`define RV_PIC_MEIPL_COUNT 12
`define RV_PIC_MEIPL_MASK 'hf
`define RV_PIC_MEIPL_OFFSET 'h0
`define RV_PIC_MEIPT_COUNT 12
`define RV_PIC_MEIPT_MASK 'h0
`define RV_PIC_MEIPT_OFFSET 'h3004
`define RV_PIC_MEIP_COUNT 4
`define RV_PIC_MEIP_MASK 'h0
`define RV_PIC_MEIP_OFFSET 'h1000
`define RV_PIC_MPICCFG_COUNT 1
`define RV_PIC_MPICCFG_MASK 'h1
`define RV_PIC_MPICCFG_OFFSET 'h3000
`define RV_PIC_OFFSET 10'hc0000
`define RV_PIC_REGION 4'hf
`define RV_PIC_SIZE 32
`define RV_PIC_TOTAL_INT 12
`define RV_PIC_TOTAL_INT_PLUS1 13
`define RV_PL2_BANK_TAGRAM_ECC_WIDTH 8
`define RV_PL2_BANK_TAGRAM_ROWS 64
`define RV_PL2_BANK_TAGRAM_WIDTH 104
`define RV_PL2_BANK_TAGRAM_WIDTH_ECC 108
`define RV_PL2_BANK_TAGRAM_WIDTH_PARITY 104
`define RV_PL2_BANK_TAG_CELL ram_64x104
`define RV_PL2_DATA_CELL ram_1024x72
`define RV_PL2_DATA_RAM_ROWS 1024
`define RV_PL2_INDEX_MSB 14
`define RV_PL2_NUM_BANKS 4
`define RV_PL2_NUM_SETS 512
`define RV_PL2_NUM_WAYS 8
`define RV_PL2_TAGRAM_ECC_64
`define RV_PL2_TAGRAM_ECC_WIDTH 8
`define RV_PL2_TAGRAM_ROWS 512
`define RV_PL2_TAGRAM_WIDTH 58
`define RV_PL2_TAGS_PER_CELL 4
`define RV_PL2_TAG_BITS 25
`define RV_PL2_TAG_CELL ram_512x58
`define RV_PL2_TAG_NUM_BANKS 8
`define RV_PLIC_BASE_ADDR 39'h68d8000000
`define RV_PLIC_IP_BASE_ADDR 39'h68dc000000
`define RV_PLIC_IP_SIZE 39'h100
`define RV_PLIC_SIZE 39'h4000000
`define RV_PMP_ENABLE
`define RV_PMP_GRAIN_MIN 4096
`define RV_PROGRAMMABLE_MISA
`define RV_RESET_CLOCK_STOP_CNTR_WIDTH 5
`define RV_RESET_VEC 'h80000000
`define RV_RET_STACK_SIZE 4
`define RV_RNMI_EXC_VEC 39'hed000000
`define RV_SB_BUS_TAG 1
`define RV_SECOND_LOAD
`define RV_SERIALIO 'hd0580000
`define RV_SHASTA_TOP shasta_wrapper
`define RV_SMODE
`define RV_STANDARD_B_EXT_EXISTS
`define RV_STANDARD_K_EXT_EXISTS
`define RV_STANDARD_ZVK_EXT_EXISTS
`define RV_STERR_ROLLBACK 0
`define RV_TARGET default
`define RV_TOP `TOP.core[0].rvtop
`define RV_TRACE_OR_AMU_EXIST
`define RV_UMODE
`define RV_UNIT_CLOCK_GATING
`define RV_UNIT_CLOCK_GATING_DEC
`define RV_UNIT_CLOCK_GATING_EXU
`define RV_UNIT_CLOCK_GATING_FPU
`define RV_UNIT_CLOCK_GATING_IFU
`define RV_UNIT_CLOCK_GATING_LSU
`define RV_UNIT_CLOCK_GATING_MMU
`define RV_UNIT_CLOCK_GATING_VEU
`define RV_UNSAFE_LOAD_STORESETS 2
`define RV_UNSAFE_LOAD_TABLE_SIZE 1024
`define RV_UNUSED_REGION0 'h0
`define RV_UNUSED_REGION1 'h10000000
`define RV_UNUSED_REGION2 'h20000000
`define RV_UNUSED_REGION3 'h30000000
`define RV_UNUSED_REGION4 'h40000000
`define RV_UNUSED_REGION5 'h50000000
`define RV_UNUSED_REGION6 'h60000000
`define RV_UNUSED_REGION7 'h70000000
`define RV_UNUSED_REGION9 'h90000000
`define RV_VEU_DEFEATURE_MAX_SEW 64
`define RV_VEU_MAX_SEW 64
`define RV_VEU_SEW_32
`define RV_VEU_SEW_64
`define RV_VIPT_ENABLE
`define SDVT_AHB 1
`define TAGE_ENTRIES_IS_2048
`define TAGE_HISTORY_SIZE 128
`define TAGE_HIST_0 2
`define TAGE_HIST_1 4
`define TAGE_HIST_10 4096
`define TAGE_HIST_11 4096
`define TAGE_HIST_12 4096
`define TAGE_HIST_13 4096
`define TAGE_HIST_14 4096
`define TAGE_HIST_2 16
`define TAGE_HIST_3 64
`define TAGE_HIST_4 128
`define TAGE_HIST_5 256
`define TAGE_HIST_6 512
`define TAGE_HIST_7 1024
`define TAGE_HIST_8 2048
`define TAGE_HIST_9 4096
`define TAGE_INDEX_WIDTH 11
`define TAGE_PRED_WIDTH 3
`define TAGE_RAM_TABLE1_FLOP 0
`define TAGE_TABLES_IS_5
`define TAGE_TAG_WIDTH 12
`define TAGE_USE_RESET_CNTR_WIDTH 18
`define TAGE_U_WIDTH 2
`define TB_BUILD_SYSREG
`define TB_CACHE_LINE_WIDTH 512
`define TB_CL_BIT_OFFSET 9
`define TB_CL_BYTE_OFFSET 6
`define TB_MMU_INDEX_TRANS
`define TB_MRAC_OVERRIDE 32'h59555555
`define TB_RV32_SYSREG_BASE_ADDR 34'hd0008000
`define TB_RV64_SYSREG_BASE_ADDR 64'h68d0008000
`define TB_SHASTA_GLOBAL_MEM_SYSTEM_MAX_CL_WIDTH_IN_BYTES 64
`define TB_SYSREG_BASE_ADDR 39'h68d0008000
`define TB_SYSREG_SIZE 39'h1000
`define TB_SYS_DCCM_OFFSET 28'h100000
`define TB_SYS_DCCM_SADR 39'h6000100000
`define TB_SYS_ICCM_OFFSET 28'h0
`define TB_SYS_ICCM_REGION 4'hc
`define TB_SYS_ICCM_SADR 39'h6000000000
`define TEC_RV_ENFLOP libenflop
`define TEC_RV_ICG clockhdr
`define TEC_RV_SYNC libsync
`define TOP tb_top
`define TOTAL_ID_SIZE 30
`define TRACE_ROUTER
`define TRC_ATDATA_BUS_WIDTH 32
`define TRC_ATID 1
`define TRC_EGRESS_FIFO_ADDR_WIDTH 4
`define TRC_IMPLICIT_RETURN_COUNTER_WIDTH 5
`define TRC_IMPLICIT_RETURN_STACK_SIZE 8
`define TRC_IMPLICIT_RETURN_STACK_WIDTH 8
`define UTLB_1G_EN
`define UTLB_NUM_WAYS 4
`define VA_SIZE 57
`define VEU_EXTERNAL_VPR
`define VPN_REQ_SIZE 47
`define VPN_SIZE 45
`define WIDE_INST_FETCH
`define TUR_AXI
`define TUR_AXI_ID_WIDTH 8
`define TUR_SOURCES 11
`define TUR_HARTS 1
`define TUR_PRIORITIES 8
`define TUR_SUPERVISOR_ENABLE
`define TUR_APLIC_M_LEVEL_CFG_BASE_ADDR 32'hd8000000
`define TUR_PLIC_BASE_ADDR 32'hd8000000
`define TOP tb_top
`define TUR_AKN_CORE_BASE_ADDR_HIGH 32'h0
`define TUR_AKN_CORE_BASE_ADDR_LOW 32'h0
`define TUR_AKN_CORE_IMSIC_MFILE_HIGH 32'h0
`define TUR_AKN_CORE_IMSIC_MFILE_LOW 32'h0
`define TUR_AKN_CORE_IMSIC_SFILE_HIGH 32'h0
`define TUR_AKN_CORE_IMSIC_SFILE_LOW 32'h0
`define TUR_AKN_CORE_IMSIC_VSFILE_HIGH 32'h0
`define TUR_AKN_CORE_IMSIC_VSFILE_LOW 32'h0
`define TUR_AKN_CORE_STRIDE_HIGH 32'h0
`define TUR_AKN_CORE_STRIDE_LOW 32'h0
`define TUR_AKN_CORE_THREAD_STRIDE 32'h0
`define TUR_APLIC_BASE_ADDR 32'hd8000000
`define TUR_APLIC_CUSTOM_AKN_BASE_ADDR 32'hd800c000
`define TUR_APLIC_M_LEVEL_IDC_BASE_ADDR 32'hd8004000
`define TUR_APLIC_S_LEVEL_CFG_BASE_ADDR 32'hd8010000
`define TUR_APLIC_S_LEVEL_IDC_BASE_ADDR 32'hd8014000
`define TUR_AXI_ADDRESS_WIDTH 32
`define TUR_AXI_SYS_ADDR_MAP {1'd0, 32'h0401_FFFF, 32'hffff_ffff}
`define TUR_AXI_SYS_ADDR_MAP_DECODE_MSB 31
`define TUR_CLINT_CSR_BASE_ADDR 32'hdc000100
`define TUR_GEILEN 0
`define TUR_IMSIC_MFILE_BASE_ADDR 32'h25000
`define TUR_IMSIC_MFILE_END_ADDR 32'h26fff
`define TUR_IMSIC_SFILE_BASE_ADDR 32'h27000
`define TUR_IMSIC_SFILE_END_ADDR 32'h28fff
`define TUR_IMSIC_VSFILE_BASE_ADDR 32'h29000
`define TUR_IMSIC_VSFILE_END_ADDR 32'h2afff
`define TUR_MSWI_BASE_ADDR 32'hdc009000
`define TUR_MTIMECMP_BASE_ADDR 32'hdc001000
`define TUR_MTIME_BASE_ADDR 32'hdc000100
`define TUR_PLIC_IP_CFG_CSR_BASE_ADDR 32'hdc000000
`define TUR_SNAPSHOT
`define TUR_SSWI_BASE_ADDR 32'hdc00d000
`define TUR_TARGETS 2
`define TUR_THREAD_PER_CORE {1'd1}, {1'd1}
`define TUR_THREAD_PER_CORE_NUM 0
`define TUR_THREAD_PER_CORE_WIDTH 0
